module xor_trigger (
    input clk,
    input rstn,
    input in, 
    output reg out
);
//在此处添加你的代码
/* always @(...)begin...
    end
*/

endmodule