module user_module (
    input clk,
    input rstn,
    input in, 
    output reg out
);
// 在此处添加您的代码
// ...

endmodule