module decimal_counter(
    input clk,
    input rstn,
    output [3:0] count
    );
    reg [3:0] q;
    assign count = q;

endmodule