module jk_ff(
    input j,
    input k,
    input clk,
    input rst,
    output q
);
reg q;
/*
always@(      )begin
    
end
*/
endmodule