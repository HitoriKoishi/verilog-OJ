
module nand3_gate(
    input a,
    input b,
    input c,
    output y
);
//在此处添加你的代码

endmodule