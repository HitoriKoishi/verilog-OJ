
module nand_gate_3(
    input a,
    input b,
    input c,
    output r
);
//在此处添加你的代码

endmodule