module user_module (
    input clk,
    input rstn,
    input in, 
    output reg out
);
// �ڴ˴�������Ĵ���
// ...

endmodule