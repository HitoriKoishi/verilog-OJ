module d_ff(
    input d,
    input clk,
    output q
    );
    reg	q; 

endmodule