
module jk_ff(
    input clk,
    input rst,
    input j,
    input k,
    output q
);
reg q;
/*
always@(      )begin
    
end
*/
endmodule