module three_vote
(
    input a,
    input b,
    input c,
    output r
);
//在此处添加你的代码

endmodule